library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;
    
package test_pkg is
    type num_array is array(natural range <>) of signed;
end package;